library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity gfp is
generic(sem_bits:natural:=3); 
port(
	modo : in std_logic
);
end entity;

architecture arch1 of gfp is
begin
end architecture;